-- Testbench de MUX 2x1bit
library IEEE;
use IEEE.std_logic_1164.all;
 
entity testbench_mux2_1bit is
end entity; 

-- Arquitetura
architecture tb of testbench_mux2_1bit is
-- Componente para DUT
component mux2_1bit is
port(
  i_sel: in std_logic;    -- entrada seletor
  i_a: in std_logic;      -- entrada a
  i_b: in std_logic;      -- entrada b
  o_q: out std_logic);    -- saída q
end component;

-- Sinais temporários
signal w_sel, w_a, w_b, w_q: std_logic;

begin
  -- Conectando os sinais no DUT
  DUT: mux2_1bit port map(
    i_sel => w_sel,
    i_a => w_a,
    i_b => w_b,
    o_q => w_q);

  process
  begin
  	w_sel <= '0';
    w_a <= '0';
    w_b <= '0';
    wait for 1 ns;
    assert(w_q='0') report "Falhou em 0/0/0" severity error;
  
    w_sel <= '1';
    w_a <= '0';
    w_b <= '0';
    wait for 1 ns;
    assert(w_q='0') report "Falhou em 1/0/0" severity error;

	  w_sel <= '0';
    w_a <= '1';
    w_b <= '0';
    wait for 1 ns;
    assert(w_q='1') report "Falhou em 0/1/0" severity error;

	  w_sel <= '0';
    w_a <= '0';
    w_b <= '1';
    wait for 1 ns;
    assert(w_q='0') report "Falhou em 0/0/1" severity error;
    
    w_sel <= '1';
    w_a <= '1';
    w_b <= '0';
    wait for 1 ns;
    assert(w_q='0') report "Falhou em 1/1/0" severity error;
    
    w_sel <= '1';
    w_a <= '0';
    w_b <= '1';
    wait for 1 ns;
    assert(w_q='1') report "Falhou em 1/0/1" severity error;
    
    w_sel <= '0';
    w_a <= '1';
    w_b <= '1';
    wait for 1 ns;
    assert(w_q='1') report "Falhou em 0/1/1" severity error;
    
    w_sel <= '1';
    w_a <= '1';
    w_b <= '1';
    wait for 1 ns;
    assert(w_q='1') report "Falhou em 1/1/1" severity error;
    
    -- Zerando entradas
    w_sel <= '0';
    w_a <= '0';
    w_b <= '0';

    assert false report "Teste feito." severity note;
    wait;
  end process;
end architecture;
